-----------------------------------------------------------------------------
--  LEON3 Demonstration design test bench
--  Copyright (C) 2004 Jiri Gaisler, Gaisler Research
------------------------------------------------------------------------------
--  This file is a part of the GRLIB VHDL IP LIBRARY
--  Copyright (C) 2003 - 2008, Gaisler Research
--  Copyright (C) 2008 - 2014, Aeroflex Gaisler
--
--  This program is free software; you can redistribute it and/or modify
--  it under the terms of the GNU General Public License as published by
--  the Free Software Foundation; either version 2 of the License, or
--  (at your option) any later version.
--
--  This program is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
--  GNU General Public License for more details.
--
--  You should have received a copy of the GNU General Public License
--  along with this program; if not, write to the Free Software
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 
------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
library gaisler;
use gaisler.libdcom.all;
use gaisler.sim.all;
library techmap;
use techmap.gencomp.all;
library micron;
use micron.components.all;
use work.debug.all;

use work.config.all;

entity testbench is
  generic (
    fabtech   : integer := CFG_FABTECH;
    memtech   : integer := CFG_MEMTECH;
    padtech   : integer := CFG_PADTECH;
    clktech   : integer := CFG_CLKTECH;
    disas     : integer := CFG_DISAS;   -- Enable disassembly to console
    dbguart   : integer := CFG_DUART;   -- Print UART on console
    pclow     : integer := CFG_PCLOW;
    clkperiod : integer := 50           -- system clock period
    );
end;

architecture behav of testbench is
  constant promfile  : string  := "prom.srec";      -- rom contents
  constant sdramfile : string  := "ram.srec";       -- sdram contents

  constant lresp    : boolean := false;
  constant ct       : integer := clkperiod/2;

  signal clk        : std_logic := '0';
  signal rst        : std_logic := '0';
  signal rstn      : std_logic;
  signal error      : std_logic;

  -- output clock
  signal clk_out    : std_ulogic;

  -- PROM flash
  signal address    : std_logic_vector(26 downto 0):=(others =>'0');
  signal data       : std_logic_vector(31 downto 0);
  signal RamCE      : std_logic;
  signal oen        : std_ulogic;
  signal writen     : std_ulogic;

  -- Debug support unit
  signal dsubre     : std_ulogic;

  -- AHB Uart
  signal dsurx      : std_ulogic;
  signal dsutx      : std_ulogic;

  -- APB Uart
  signal rxd1       : std_ulogic;
  signal txd1       : std_ulogic;

  -- Output signals for LEDs
  signal led       : std_logic_vector(1 downto 0);
  signal gpio      : std_logic_vector(7 downto 0);

  -- Output signals for LEDs
  signal triggerout : std_logic_vector(3 downto 0);
  signal alarmout   : std_ulogic;
  signal alarmin   : std_ulogic;
  signal clkout : std_ulogic;
  signal extsave     : std_ulogic;

begin
  -- clock and reset
  clk        <= not clk after ct * 1 ns;
  rst        <= '1', '0' after 100 ns;
  rstn       <= rst;
  dsubre     <= '0';
  rxd1      <= 'H';
  
  d3 : entity work.leon3mp
    --generic map (fabtech, memtech, padtech, clktech)
    port map (
      clk     => clk,
      btnCpuResetn => rstn,
      
     -- output signals for led
      led => led,
      gpio => gpio,
      errorn => error,
      
      -- PROM
     --address   => address(22 downto 0),
     --data      => data(31 downto 16),
     --
     --RamOE     => oen,
     --RamWE     => writen,
     --RamCE     => RamCE,
  
      -- APB Uart
      rxd1 => rxd1,
      txd1 => txd1,

      -- AHB Uart
      RsRx     => dsurx,
      RsTx     => dsutx,
      
      alarmin => alarmin,
      clkout => clkout,
      triggerout =>  triggerout,
      alarmout => alarmout,
      extsave => extsave

      );

  --sram0 : sram
    --generic map (index => 4, abits => 24, fname => sdramfile)
    --port map (address(23 downto 0), data(31 downto 24), RamCE, writen, oen);

  --sram1 : sram
    --generic map (index => 5, abits => 24, fname => sdramfile)
    --port map (address(23 downto 0), data(23 downto 16), RamCE, writen, oen);

     
  extsave <= 'L';

  iuerr : process
  begin
    wait for 5 us;
    assert (to_X01(error) = '1')
      report "*** IU in error mode, simulation halted ***"
      severity failure;
  end process;

  data <= buskeep(data) after 5 ns;

 end;
